module top(in_data, out_data);
  bit [1:0] _00_;
  bit [1:0] _01_;
  bit _02_;
  bit _03_;
  bit _04_;
  bit _05_;
  bit [1:0] _06_;
  bit [1:0] _07_;
  bit _08_;
  bit _09_;
  bit _10_;
  bit celloutsig_0z;
  bit [1:0] celloutsig_1z;
  bit [1:0] celloutsig_2z;
  bit celloutsig_3z;
  input [95:0] in_data;
  bit [95:0] in_data;
  output [95:0] out_data;
  bit [95:0] out_data;
  assign celloutsig_1z = _01_ * _00_;
  assign celloutsig_2z = _05_ ? _06_ : _07_;
  assign celloutsig_3z = _02_ ? _03_ : _04_;
  assign celloutsig_0z = _09_ | _08_;
  assign _09_ = in_data[21];
  assign _08_ = in_data[51];
  assign _01_[0] = celloutsig_0z;
  assign _01_[1] = celloutsig_0z;
  assign _00_[0] = celloutsig_0z;
  assign _00_[1] = celloutsig_0z;
  assign _07_[0] = celloutsig_0z;
  assign _07_[1] = celloutsig_1z[0];
  assign _06_ = in_data[43:42];
  assign _05_ = celloutsig_1z[0];
  assign _04_ = celloutsig_2z[1];
  assign _03_ = celloutsig_2z[0];
  assign _02_ = in_data[43];
  assign _10_ = in_data[92];
  assign out_data[32] = celloutsig_3z;
endmodule
